build_base_covmodel_tree();
