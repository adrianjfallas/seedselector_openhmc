`include "seed_selector/cov_tree_defs_and_methods.sv"

function void build_base_covmodel_tree();

	$display("SEED_SELECTOR: First test run, no coverage tree yet.");

endfunction
