`include "seed_selector/cov_tree_defs_and_methods.sv"

function int build_base_covmodel_tree(int influence_param_1);

	$display("SEED_SELECTOR: First test run, no coverage tree yet.");

endfunction
